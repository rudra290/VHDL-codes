-- A DUT entity is used to wrap your design.
--  This example shows how you can do this for the
--  Full-adder.

library ieee;
use ieee.std_logic_1164.all;

entity DUT is
   port(input_vector: in std_logic_vector(8 downto 0);
       	output_vector: out std_logic_vector(7 downto 0));
end entity;

architecture DutWrap of DUT is
	-- Instantiate your own top Module component in place of ALU_1
	
component Quiz is
port( A : in std_logic_vector(7 downto 0);
		M : in std_logic;
		Y : out std_logic_vector(7 downto 0)
	 );
end component;

begin

   -- input/output vector element ordering is critical,
   -- and must match the ordering in the trace file!
   dut_instance: Quiz port map (M => input_vector(8), A(7 downto 0) => input_vector(7 downto 0),
										  y(7 downto 0) => output_vector(7 downto 0));

end DutWrap;

